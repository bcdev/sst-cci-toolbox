netcdf aai_20101224 {
dimensions:
	nx = 288 ;
	ny = 180 ;
variables:
	float lon(nx) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
	float lat(ny) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
	float aerosol_absorbing_index(ny, nx) ;
		aerosol_absorbing_index:long_name = "Aerosol: Absorbing Aerosol Index" ;
		aerosol_absorbing_index:units = "percent" ;
		aerosol_absorbing_index:_FillValue = -32768.f ;

// global attributes:
		:title = "Global Aerosol - Absorbing Aerosol Index" ;
		:institution = "University of Leicester" ;
		:contact = "Christopher Whyte (ce101@le.ac.uk)" ;
		:creation_date = "Tue May 17 10:32:00 2011" ;
		:callsign = "GOME-2" ;
}
