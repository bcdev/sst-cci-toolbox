netcdf l4 {
dimensions:
    lon = 7200 ;
    lat = 3600 ;
    time = 1 ;
    bnds = 2 ;
variables:
    float lat(lat) ;
        lat:units = "degrees_north" ;
        lat:long_name = "Latitude coordinates" ;
        lat:standard_name = "latitude" ;
        lat:valid_min = -90.0f ;
        lat:valid_max = 90.0f ;
        lat:reference_datum = "geographical coordinates, WGS84 projection" ;
        lat:axis = "Y" ;
        lat:bounds = "lat_bnds" ;
    float lat_bnds(lat, bnds) ;
        lat_bnds:units = "degrees_north" ;
        lat_bnds:long_name = "Latitude cell boundaries" ;
        lat_bnds:valid_min = -90.0f ;
        lat_bnds:valid_max = 90.0f ;
        lat_bnds:reference_datum = "geographical coordinates, WGS84 projection" ;
        lat_bnds:comment = "Contains the northern and southern boundaries of the grid cells";
    float lon(lon) ;
        lon:units = "degrees_east" ;
        lon:long_name = "Longitude coordinates" ;
        lon:standard_name = "longitude" ;
        lon:valid_min = -180.0f ;
        lon:valid_max = 180.0f ;
        lon:reference_datum = "geographical coordinates, WGS84 projection" ;
        lat:axis = "X" ;
        lat:bounds = "lon_bnds" ;
    float lon_bnds(lon, bnds) ;
        lon_bnds:units = "degrees_east" ;
        lon_bnds:long_name = "Longitude cell boundaries" ;
        lon_bnds:valid_min = -90.0f ;
        lon_bnds:valid_max = 90.0f ;
        lon_bnds:reference_datum = "geographical coordinates, WGS84 projection" ;
        lon_bnds:comment = "Contains the western and eastern boundaries of the grid cells";
    int time(time) ;
        time:units = "seconds since 1981-01-01 00:00:00" ;
        time:long_name = "reference time of sst file" ;
        time:standard_name = "time" ;
        time:calendar = "gregorian" ;
        time:axis = "T" ;
        time:bounds = "time_bnds" ;
    float time_bnds(time, bnds) ;
        time_bnds:units = "seconds since 1981-01-01 00:00:00" ;
        time_bnds:long_name = "Time cell boundaries" ;
        time_bnds:calendar = "gregorian" ;
        time_bnds:comment = "Contains the start and end times for the time period the data represent";
    short analysed_sst(time, lat, lon) ;
        analysed_sst:_FillValue = -32768s ;
        analysed_sst:units = "kelvin" ;
        analysed_sst:scale_factor = 0.01f ;
        analysed_sst:add_offset = 273.15f ;
        analysed_sst:long_name = "analysed sea surface temperature" ;
        analysed_sst:valid_min = -300s;
        analysed_sst:valid_max = 4500;
        analysed_sst:standard_name = "sea_surface_foundation_temperature" ;
        analysed_sst:source = "TBD" ;
        analysed_sst:depth = "20 cm" ;
    short analysis_error(time, lat, lon) ;
        analysis_error:_FillValue = -32768s ;
        analysis_error:units = "kelvin" ;
        analysis_error:scale_factor = 0.01f ;
        analysis_error:add_offset = 0.0f ;
        analysis_error:long_name = "Estimated error standard deviation of analysed_sst" ;
        analysis_error:valid_min = 0s ;
        analysis_error:valid_max = 32767s ;
        analysis_error:standard_name = "sea_surface_foundation_temperature_standard_error" ;
    byte sea_ice_fraction(time, lat, lon) ;
        sea_ice_fraction:_FillValue = -128b ;
        sea_ice_fraction:units = "1" ;
        sea_ice_fraction:scale_factor = 0.01f ;
        sea_ice_fraction:add_offset = 0.0f ;
        sea_ice_fraction:long_name = "Sea ice area fraction" ;
        sea_ice_fraction:valid_min = 0b ;
        sea_ice_fraction:valid_max = 100b ;
        analysis_error:standard_name = "sea_ice_area_fraction" ;
        sea_ice_fraction:comment = "Component of uncertainty that is correlated over synoptic scales; can be combined with other uncertainty estimates to form a total uncertainty" ;
        sea_ice_fraction:source = "EUMETSAT_OSI_SAF-ICE-v<TBC>" ;
    byte mask(time, lat, lon) ;
        mask:long_name = "sea/land/lake/ice field composite mask" ;
        mask:comment = "b0: 1=grid cell is open sea water b1: 1=land is present in this grid cell b2: 1=lake surface is present in this grid cell b3: 1=sea ice is present in this grid cell b4-b7: reserved for future grid mask data" ;
        mask:flag_meanings = "sea land lake ice" ;
        mask:flag_masks = 1b, 2b, 4, 8b ;

// global attributes:
        :Conventions = "CF-1.4" ;
        :title = "ESA SST CCI OSTIA L4 product" ;
        :summary = "OSTIA L4 product from the ESA SST CCI project, produced using <algorithm name>" ;
        :references = "TBD" ;
        :institution = "ESACCI" ;
        :history = "" ;
        :license = "GHRSST protocol describes data use as free and open" ;
        :id = "TBD" ;
        :naming_authority = "org.ghrsst" ;
        :product_version = "TBD" ;
        :uuid = "TBD" ;
        :gds_version_id = "2.0" ;
        :netcdf_version_id = "4.1.3" ;
        :date_created = "20120131T120000Z" ;
        :file_quality_level = 0 ;
        :spatial_resolution = "1 km" ;
        :start_time = "20120131070000Z" ;
        :time_coverage_start = "20120131070000Z" ;
        :stop_time = "20120131083000Z" ;
        :source = "AATSR-ESA-L1-v2.0" ;
        :platform = "" ;
        :sensor = "OSTIA (analysis)" ;
        :metadata_conventions = "Unidata Dataset Discovery v1.0" ;
        :metadata_link = "TBD" ;
        :keywords = "Oceans > Ocean > Temperature > Sea Surface Temperature" ;
        :keywords_vocabulary = "NASA Global Change Master Directory (GCMD) Science Keywords" ;
        :standard_name_vocabulary = "NetCDF Climate and Forecast (CF) Metadata Convention" ;
        :geospatial_lat_units = "degrees_north" ;
        :geospatial_lat_resolution = 0.05f ;
        :geospatial_lon_units = "degrees_east" ;
        :geospatial_lon_resolution = 0.05f ;
        :acknowledgment = "Funded by ESA" ;
        :creator_name = "ESA SST CCI" ;
        :creator_email = "science.lead er@esa-sst- cci.org" ;
        :creator_url = "http://www.es a-sst-cci.org/" ;
        :project = "European Space Agency Sea Surface Temperature Climate Change Initiative" ;
        :publisher_name = "The GHRSST Project Office" ;
        :publisher_email = "ghrsst- po@nceo.ac.uk" ;
        :publisher_url = "http://www.g hrsst.org" ;
        :comment = "These data were produced at <institution> as part of the ESA SST CCI project" ;
        :northernmost_latitude = 90.0f ;
        :southernmost_latitude = -90.0f ;
        :easternmost_longitude = 180.0f ;
        :westernmost_longitude = -180.0f ;
        :processing_level = "L4" ;
        :cdm_data_type = "grid" ;
}