netcdf 20100701000000-ESACCI-L4_GHRSST-SSTdepth-OSTIA-LT-v02.0-fv01.0 {
dimensions:
	lon = 7200 ;
	lat = 3600 ;
	bnds = 2 ;
	time = UNLIMITED ; // (0 currently)
variables:
	float lat(lat) ;
		lat:units = "degrees_north" ;
		lat:long_name = "Latitude" ;
		lat:standard_name = "latitude" ;
		lat:valid_min = -90.f ;
		lat:valid_max = 90.f ;
		lat:reference_datum = "geographical coordinates, WGS84 projection" ;
		lat:axis = "Y" ;
		lat:bounds = "lat_bnds" ;
	float lat_bnds(lat, bnds) ;
		lat_bnds:units = "degrees_north" ;
		lat_bnds:long_name = "Latitude cell boundaries" ;
		lat_bnds:valid_min = -90.f ;
		lat_bnds:valid_max = 90.f ;
		lat_bnds:comment = "Contains the northern and southern boundaries of the grid cells." ;
		lat_bnds:reference_datum = "geographical coordinates, WGS84 projection" ;
	float lon(lon) ;
		lon:units = "degrees_east" ;
		lon:long_name = "Longitude" ;
		lon:standard_name = "longitude" ;
		lon:valid_min = -180.f ;
		lon:valid_max = 180.f ;
		lon:reference_datum = "geographical coordinates, WGS84 projection" ;
		lon:axis = "X" ;
		lon:bounds = "lon_bnds" ;
	float lon_bnds(lon, bnds) ;
		lon_bnds:units = "degrees_east" ;
		lon_bnds:long_name = "Longitude cell boundaries" ;
		lon_bnds:valid_min = -180.f ;
		lon_bnds:valid_max = 180.f ;
		lon_bnds:comment = "Contains the eastern and western boundaries of the grid cells." ;
		lon_bnds:reference_datum = "geographical coordinates, WGS84 projection" ;
	int time(time) ;
		time:units = "seconds since 1981-01-01 00:00:00" ;
		time:long_name = "reference time of sst file" ;
		time:standard_name = "time" ;
		time:axis = "T" ;
		time:calendar = "gregorian" ;
		time:bounds = "time_bnds" ;
	float time_bnds(time, bnds) ;
		time_bnds:units = "seconds since 1981-01-01 00:00:00" ;
		time_bnds:long_name = "Time cell boundaries" ;
		time_bnds:comment = "Contains the start and end times for the time period the data represent" ;
	short analysed_sst(time, lat, lon) ;
		analysed_sst:_FillValue = -32768s ;
		analysed_sst:units = "kelvin" ;
		analysed_sst:scale_factor = 0.01f ;
		analysed_sst:add_offset = 273.15f ;
		analysed_sst:long_name = "analysed sea surface temperature" ;
		analysed_sst:valid_min = -300s ;
		analysed_sst:valid_max = 4500s ;
		analysed_sst:standard_name = "sea_water_temperature" ;
		analysed_sst:source = "AATSR-ESACCI-L3U-LT-v01.0, AVHRR19_G- ESACCI-L2P-LT-v01.0" ;
		analysed_sst:depth = "20 cm" ;
	short analysis_error(time, lat, lon) ;
		analysis_error:_FillValue = -32768s ;
		analysis_error:units = "kelvin" ;
		analysis_error:scale_factor = 0.01f ;
		analysis_error:add_offset = 0.f ;
		analysis_error:long_name = "estimated error standard deviation of analysed_sst" ;
		analysis_error:valid_min = 0s ;
		analysis_error:valid_max = 32767s ;
		analysis_error:standard_name = "sea_water_temperature standard_error" ;
	byte sea_ice_fraction(time, lat, lon) ;
		sea_ice_fraction:_FillValue = -128b ;
		sea_ice_fraction:units = "1" ;
		sea_ice_fraction:scale_factor = 0.01f ;
		sea_ice_fraction:add_offset = 0.f ;
		sea_ice_fraction:long_name = "sea ice area fraction" ;
		sea_ice_fraction:valid_min = 0s ;
		sea_ice_fraction:valid_max = 100s ;
		sea_ice_fraction:standard_name = "sea_ice_area_fraction" ;
		sea_ice_fraction:source = "EUMETSAT_OSISAF-ICE-v1.1" ;
	byte mask(time, lat, lon) ;
		mask:long_name = "sea/land/lake/ice field composite mask" ;
		mask:comment = "b0: 1=grid cell is open sea water b1: 1=land is present in this grid cell b2: 1=lake surface is present in this grid cell b3: 1=sea ice is present in this grid cell b4-b7: reserved for future grid mask data" ;
		mask:flag_meanings = "sea land lake ice" ;
		mask:flag_values = 1b, 2b, 4b, 8b ;
data:
    lat = ${LAT} ;
    lon = ${LON} ;

// global attributes:
		:Conventions = "CF-1.5, Unidata Observation Dataset v1.0" ;
		:title = "ESA SST CCI OSTIA L4 product" ;
		:summary = "OSTIA L4 product from the ESA SST CCI project, produced using <algorithm name>." ;
		:references = "Insert published or web-based references that\n",
			"describe the data or methods used to produce them" ;
		:institution = "ESACCI" ;
		:history = "SST CCI processor XXX.YY" ;
		:licence = "TBC" ;
		:id = "OSTIA-ESACCI-L4-v<Version Number>" ;
		:naming_authority = "org.ghrsst" ;
		:product_version = "1.0" ;
		:uuid = "D7A88FA8-7421-4039-807C-B551D638EDC6" ;
		:tracking_id = "D7A88FA8-7421-4039-807C-B551D638EDC6" ;
		:gds_version_id = "2.0" ;
		:netcdf_version_id = "4.1.1" ;
		:date_created = "20110616T152836Z" ;
		:file_quality_level = 3 ;
		:spatial_resolution = "1.1km at nadir" ;
		:start_time = "20100701T000000Z" ;
		:time_coverage_start = "20100701T000000Z" ;
		:stop_time = "20100701T235959Z" ;
		:time_coverage_end = "20100701T235959Z" ;
		:time_coverage_duration = "P1D" ;
		:time_coverage_resolution = "P1D" ;
		:source = "AATSR-ESACCI-L3U-v1.0, AVHRR-ESACCI-L2P-v1.0, EUMETSAT_OSISAF-ICE-v1.1" ;
		:platform = "Envisat, NOAA-<X>" ;
		:sensor = "AATSR" ;
		:metadata_conventions = "Unidata Dataset Discovery v1.0" ;
		:metadata_link = "http://www.esa-cci.org" ;
		:keywords = "Oceans > Ocean Temperature > Sea Surface Temperature" ;
		:keywords_vocabulary = "NASA Global Change Master Directory (GCMD) Science Keywords" ;
		:standard_name_vocabulary = "NetCDF Climate and Forecast (CF) Metadata Convention" ;
		:geospatial_lat_units = "degrees_north" ;
		:geospatial_lat_resolution = "0.05" ;
		:geospatial_lon_units = "degrees_east" ;
		:geospatial_lon_resolution = "0.05" ;
		:geospatial_vertical_min = -0.2f ;
		:geospatial_vertical_max = -0.2f ;
		:acknowledgment = "Funded by ESA" ;
		:creator_name = "ESA SST CCI" ;
		:creator_email = "science.leader@esa-sst-cci.org" ;
		:creator_url = "http://www.esa-sst-cci.org" ;
		:creator_processing_institution = "These data were produced at the Met Office as part of the ESA SST CCI project." ;
		:project = "European Space Agency Sea Surface Temperature Climate Change Initiative" ;
		:publisher_name = "ESACCI" ;
		:publisher_url = "http://www.esa-sst-cci.org" ;
		:publisher_email = "science.leader@esa-SST-cci.org" ;
		:comment = "" ;
		:northernmost_latitude = 90.f ;
		:southernmost_latitude = -90.f ;
		:easternmost_longitude = -180.f ;
		:westernmost_longitude = 180.f ;
		:geospatial_lat_max = 90.f ;
		:geospatial_lat_min = -90.f ;
		:geospatial_lon_max = -180.f ;
		:geospatial_lon_min = 180.f ;
		:processing_level = "L4" ;
		:cdm_data_type = "grid" ;
}
