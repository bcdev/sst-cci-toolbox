netcdf 20100701000000-ESACCI-L2P_GHRSST-SSTskin-AATSR-DM-v02.0-fv01.0 {
dimensions:
	ni = 512 ;
	nj = 28000 ;
	time = 1 ;
variables:
	float lat(nj, ni) ;
		lat:units = "degrees_north" ;
		lat:long_name = "Latitude coordinates" ;
		lat:standard_name = "latitude" ;
		lat:valid_min = -90.f ;
		lat:valid_max = 90.f ;
		lat:reference_datum = "geographical coordinates, WGS84 projection" ;
	float lon(nj, ni) ;
		lon:units = "degrees_east" ;
		lon:long_name = "Longitude coordinates" ;
		lon:standard_name = "longitude" ;
		lon:valid_min = -180.f ;
		lon:valid_max = 180.f ;
		lon:reference_datum = "geographical coordinates, WGS84 projection" ;
	int time(time) ;
		time:units = "seconds since 1981-01-01 00:00:00" ;
		time:long_name = "reference time of sst file" ;
		time:standard_name = "time" ;
		time:calendar = "gregorian" ;
	short sea_surface_temperature(time, nj, ni) ;
		sea_surface_temperature:_FillValue = -32768s ;
		sea_surface_temperature:units = "kelvin" ;
		sea_surface_temperature:scale_factor = 0.01f ;
		sea_surface_temperature:add_offset = 273.15f ;
		sea_surface_temperature:long_name = "sea surface skin temperature" ;
		sea_surface_temperature:valid_min = -200s ;
		sea_surface_temperature:valid_max = 5000s ;
		sea_surface_temperature:standard_name = "sea_surface_skin_temperature" ;
		sea_surface_temperature:comment = "Temperature of the skin of the ocean; total uncertainty = sqrt(large_scale_correlated_uncertainty^2 + synoptically_correlated_uncert ainty^2 + uncorrelated_uncertainty^2)" ;
		sea_surface_temperature:source = "AATSR-ESA-L1-v2.0" ;
		sea_surface_temperature:references = "Insert published or web-based references that describe the data or methods used to produce them" ;
		sea_surface_temperature:depth = "10 micrometres" ;
		sea_surface_temperature:coordinates = "lon lat" ;
	short sst_dtime(time, nj, ni) ;
		sst_dtime:_FillValue = -32768s ;
		sst_dtime:units = "seconds" ;
		sst_dtime:scale_factor = 1.f ;
		sst_dtime:add_offset = 0.f ;
		sst_dtime:long_name = "time difference from reference time" ;
		sst_dtime:valid_min = -32767s ;
		sst_dtime:valid_max = 32767s ;
		sst_dtime:comment = "time plus sst_dtime gives seconds after 1981-01-01 00:00:00" ;
		sst_dtime:coordinates = "lon lat" ;
	byte sses_bias(time, nj, ni) ;
		sses_bias:_FillValue = -128b ;
		sses_bias:units = "kelvin" ;
		sses_bias:scale_factor = 0.01f ;
		sses_bias:add_offset = 0.f ;
		sses_bias:long_name = "SSES bias estimate" ;
		sses_bias:valid_min = -127b ;
		sses_bias:valid_max = 127b ;
		sses_bias:comment = "Populated with zeroes" ;
		sses_bias:coordinates = "lon lat" ;
	byte sses_standard_deviation(time, nj, ni) ;
		sses_standard_deviation:_FillValue = -128b ;
		sses_standard_deviation:units = "kelvin" ;
		sses_standard_deviation:scale_factor = 0.01f ;
		sses_standard_deviation:add_offset = 0.f ;
		sses_standard_deviation:long_name = "SSES standard deviation" ;
		sses_standard_deviation:valid_min = -127b ;
		sses_standard_deviation:valid_max = 127b ;
		sses_standard_deviation:comment = "Total uncertainty in each sea_surface_temperature data point" ;
		sses_standard_deviation:coordinates = "lon lat" ;
	short l2p_flags(time, nj, ni) ;
		l2p_flags:long_name = "L2P flags" ;
		l2p_flags:comment = "These flags are important to properly use the data" ;
		l2p_flags:coordinates = "lon lat" ;
		l2p_flags:flag_meanings = "microwave land ice lake river spare views channels" ;
		l2p_flags:flag_masks = 1s, 2s, 4s, 8s, 16s, 32s, 64s, 128s ;
	byte quality_level(time, nj, ni) ;
		quality_level:long_name = "quality level of SST pixel" ;
		quality_level:comment = "These are overall quality indicators and are those used for all GHRSST SSTs" ;
		quality_level:coordinates = "lon lat" ;
		quality_level:flag_meanings = "no_data bad_data worst_quality low_quality acceptable_quality best_quality" ;
		quality_level:flag_values = 0b, 1b, 2b, 3b, 4b, 5b ;
	byte wind_speed(time, nj, ni) ;
		wind_speed:_FillValue = -128b ;
		wind_speed:units = "m s-1" ;
		wind_speed:scale_factor = 0.1f ;
		wind_speed:add_offset = 12.7f ;
		wind_speed:long_name = "10m wind speed" ;
		wind_speed:valid_min = -127b ;
		wind_speed:valid_max = 127b ;
		wind_speed:standard_name = "wind_speed" ;
		wind_speed:comment = "Wind speeds sourced from ECMWF ERA Interim reanalysis; wind speeds greater than 25.4 m/s are set to 25.4" ;
		wind_speed:source = "ERA_INTERIM-ECMWF-WSP-v1.0" ;
		wind_speed:references = "Insert published or web-based references that describe the data or methods used to produce them" ;
		wind_speed:coordinates = "lon lat" ;
		wind_speed:height = "10 m" ;
		wind_speed:time_offset = 1.f ;
	short sea_surface_temperature_depth(time, nj, ni) ;
		sea_surface_temperature_depth:_FillValue = -32768s ;
		sea_surface_temperature_depth:units = "kelvin" ;
		sea_surface_temperature_depth:scale_factor = 0.01f ;
		sea_surface_temperature_depth:add_offset = 273.15f ;
		sea_surface_temperature_depth:long_name = "sea surface temperature at 0.2 m" ;
		sea_surface_temperature_depth:valid_min = -200s ;
		sea_surface_temperature_depth:valid_max = 5000s ;
		sea_surface_temperature_depth:standard_name = "sea_water_temperature" ;
		sea_surface_temperature_depth:comment = "Temperature of the ocean at 20 cm depth; total uncertainty = sqrt(large_scale_correlated_uncertainty^2 + synoptically_correlated_uncertainty^2 + uncorrelated_uncertainty^2 + adjustment_uncertainty^2)" ;
		sea_surface_temperature_depth:source = "AATSR-ESA-L1-v2.0" ;
		sea_surface_temperature_depth:references = "Insert published or web-based references that describe the data or methods used to produce them" ;
		sea_surface_temperature_depth:depth = "0.2 metre" ;
		sea_surface_temperature_depth:coordinates = "lon lat" ;
	short large_scale_correlated_uncertainty(time, nj, ni) ;
		large_scale_correlated_uncertainty:_FillValue = -32768s ;
		large_scale_correlated_uncertainty:units = "kelvin" ;
		large_scale_correlated_uncertainty:scale_factor = 0.01f ;
		large_scale_correlated_uncertainty:add_offset = 0.f ;
		large_scale_correlated_uncertainty:long_name = "Uncertainty from errors likely to be correlated over large scales" ;
		large_scale_correlated_uncertainty:valid_min = 0s ;
		large_scale_correlated_uncertainty:valid_max = 5000s ;
		large_scale_correlated_uncertainty:comment = "Component of uncertainty that is correlated over large scales; can be combined with other uncertainty estimates to form a total uncertainty" ;
		large_scale_correlated_uncertainty:references = "Insert published or web-based references that describe the data or methods used to produce them" ;
		large_scale_correlated_uncertainty:coordinates = "lon lat" ;
	short synoptically_correlated_uncertainty(time, nj, ni) ;
		synoptically_correlated_uncertainty:_FillValue = -32768s ;
		synoptically_correlated_uncertainty:units = "kelvin" ;
		synoptically_correlated_uncertainty:scale_factor = 0.01f ;
		synoptically_correlated_uncertainty:add_offset = 0.f ;
		synoptically_correlated_uncertainty:long_name = "Uncertainty from errors likely to be correlated over synoptic scales" ;
		synoptically_correlated_uncertainty:valid_min = 0s ;
		synoptically_correlated_uncertainty:valid_max = 5000s ;
		synoptically_correlated_uncertainty:comment = "Component of uncertainty that is correlated over synoptic scales; can be combined with other uncertainty estimates to form a total uncertainty" ;
		synoptically_correlated_uncertainty:references = "Insert published or web-based references that describe the data or methods used to produce them" ;
		synoptically_correlated_uncertainty:coordinates = "lon lat" ;
		synoptically_correlated_uncertainty:correlation_length_scale = "100 km" ;
		synoptically_correlated_uncertainty:correlation_time_scale = "1 day" ;
	short uncorrelated_uncertainty(time, nj, ni) ;
		uncorrelated_uncertainty:_FillValue = -32768s ;
		uncorrelated_uncertainty:units = "kelvin" ;
		uncorrelated_uncertainty:scale_factor = 0.01f ;
		uncorrelated_uncertainty:add_offset = 0.f ;
		uncorrelated_uncertainty:long_name = "Uncertainty from errors likely to be uncorrelated between SSTs" ;
		uncorrelated_uncertainty:valid_min = 0s ;
		uncorrelated_uncertainty:valid_max = 5000s ;
		uncorrelated_uncertainty:comment = "Component of uncertainty that is uncorrelated between SSTs; can be combined with other uncertainty estimates to form a total uncertainty" ;
		uncorrelated_uncertainty:references = "Insert published or web-based references that describe the data or methods used to produce them" ;
		uncorrelated_uncertainty:coordinates = "lon lat" ;
	short adjustment_uncertainty(time, nj, ni) ;
		adjustment_uncertainty:_FillValue = -32768s ;
		adjustment_uncertainty:units = "kelvin" ;
		adjustment_uncertainty:scale_factor = 0.01f ;
		adjustment_uncertainty:add_offset = 0.f ;
		adjustment_uncertainty:long_name = "Time and depth adjustment uncertainty" ;
		adjustment_uncertainty:valid_min = 0s ;
		adjustment_uncertainty:valid_max = 5000s ;
		adjustment_uncertainty:comment = "Adjustment uncertainty; can be combined with other uncertainty estimates to form a total uncertainty" ;
		adjustment_uncertainty:references = "Insert published or web-based references that describe the data or methods used to produce them" ;
		adjustment_uncertainty:coordinates = "lon lat" ;
		adjustment_uncertainty:correlation_length_scale = "100 km" ;
		adjustment_uncertainty:correlation_time_scale = "1 day" ;

// global attributes:
		:Conventions = "CF-1.5" ;
		:title = "ESA SST CCI AATSR L2P product" ;
		:summary = "AATSR L2P product from the ESA SST CCI project, produced using <algorithm name>." ;
		:references = "Insert published or web-based references that describe the data or methods used to produce them" ;
		:institution = "ESACCI" ;
		:history = "SST CCI processor XXX.YY" ;
		:licence = "TBC" ;
		:id = "AATSR-ESACCI-L2P-v<Version Number>" ;
		:naming_authority = "org.ghrsst" ;
		:product_version = "1.0" ;
		:uuid = "D7A88FA8-7421-4039-807C-B551D638EDC6" ;
		:tracking_id = "D7A88FA8-7421-4039-807C-B551D638EDC6" ;
		:gds_version_id = "2.0" ;
		:netcdf_version_id = "4.1.3" ;
		:date_created = "20110616T152207Z" ;
		:file_quality_level = 3 ;
		:spatial_resolution = "1.1km at nadir" ;
		:start_time = "20100701T000000Z" ;
		:time_coverage_start = "20100701T000000Z" ;
		:stop_time = "20100701T013000Z" ;
		:time_coverage_end = "20100701T013000Z" ;
		:time_coverage_duration = "PT1H30M" ;
		:time_coverage_resolution = "PT1S" ;
		:source = "AATSR-ESA-L1-v2.0, ERA_INTERIM-ECMWF-WSP-v1.0" ;
		:platform = "Envisat" ;
		:sensor = "AATSR" ;
		:metadata_conventions = "Unidata Dataset Discovery v1.0" ;
		:metadata_link = "http://www.esa-cci.org" ;
		:keywords = "Oceans > Ocean Temperature > Sea Surface Temperature" ;
		:keywords_vocabulary = "NASA Global Change Master Directory (GCMD) Science Keywords" ;
		:standard_name_vocabulary = "NetCDF Climate and Forecast (CF) Metadata Convention" ;
		:geospatial_lat_units = "degrees_north" ;
		:geospatial_lat_resolution = "0.009" ;
		:geospatial_lon_units = "degrees_east" ;
		:geospatial_lon_resolution = "0.009" ;
		:geospatial_vertical_min = -0.2f ;
		:geospatial_vertical_max = -1.e-05f ;
		:acknowledgment = "Funded by ESA" ;
		:creator_name = "ESACCI" ;
		:creator_email = "science.leader@esa-sst-cci.org" ;
		:creator_url = "http://www.esa-sst-cci.org" ;
		:creator_processing_institution = "University of Edinburgh" ;
		:project = "Climate Change Initiative - European Space Agency" ;
		:publisher_name = "ESACCI" ;
		:publisher_url = "http://www.esa-sst-cci.org" ;
		:publisher_email = "science.leader@esa-SST-cci.org" ;
		:comment = "See the comment attributes to the sea_surface_temperature and sea_surface_temperature_depth variables for information about uncertainty estimates." ;
		:northernmost_latitude = 90.f ;
		:southernmost_latitude = -90.f ;
		:easternmost_longitude = -180.f ;
		:westernmost_longitude = 180.f ;
		:geospatial_lat_max = 90.f ;
		:geospatial_lat_min = -90.f ;
		:geospatial_lon_max = -180.f ;
		:geospatial_lon_min = 180.f ;
		:processing_level = "L2P" ;
		:cdm_data_type = "swath" ;
data:
    lat = ${LAT} ;
    lon = ${LON} ;
}
