netcdf NSS.GHRR.NK.D10152.S1852.E2020.B6265657.WI.MMM {
dimensions:
	ni = 25 ;
	nj = 31 ;
	charlen = 50 ;
	matchup = UNLIMITED ; // (45 currently)
variables:
	int matchup_id(matchup) ;
	int matchup_elem(matchup) ;
		matchup_elem:orientation = "elem (1) is L1B file element (matchup_elem - 12)" ;
	int matchup_line(matchup) ;
		matchup_line:orientation = "line (1) is L1B file line (matchup_line - 15)" ;
	byte bad_data(matchup, nj, ni) ;
		bad_data:values = "0=good but individual channels may be bad; 1=bad" ;
	byte cloud_flag(matchup, nj, ni) ;
		cloud_flag:values = "bit 2:0=cloud mask valid, 1=cloud mask not valid; bits 1-0: CLAVR-x bayesian cloud mask 0=clear, 1=probably clear, 2=probably cloud, 3=cloud" ;
		cloud_flag:missing_value = 7 ;
	byte cloud_prob(matchup, nj, ni) ;
		cloud_prob:values = "CLAVR-x bayesian cloud prob, 0.0:1.0 scaled to -127:127" ;
		cloud_prob:missing_value = -128 ;
	char avhrr_name(matchup, charlen) ;
	char l1b_filename(matchup, charlen) ;
	float ict_temp(matchup, nj) ;
		ict_temp:units = "K" ;
		ict_temp:missing_value = -1.e+030f ;
	float reflec_to_rad_1(matchup) ;
		reflec_to_rad_1:units = "-" ;
		reflec_to_rad_1:missing_value = -1.e+030f ;
	float reflec_to_rad_2(matchup) ;
		reflec_to_rad_2:units = "-" ;
		reflec_to_rad_2:missing_value = -1.e+030f ;
	float reflec_to_rad_3a(matchup) ;
		reflec_to_rad_3a:units = "-" ;
		reflec_to_rad_3a:missing_value = -1.e+030f ;
	int time_year(matchup, nj) ;
		time_year:units = "year" ;
		time_year:missing_value = -32768 ;
	int time_day_num(matchup, nj) ;
		time_day_num:units = "day" ;
		time_day_num:missing_value = -32768 ;
	int time_utc_msecs(matchup, nj) ;
		time_utc_msecs:units = "msec" ;
		time_utc_msecs:missing_value = -32768 ;
	float longitude(matchup, nj, ni) ;
		longitude:units = "deg" ;
		longitude:missing_value = -1.e+030f ;
	float latitude(matchup, nj, ni) ;
		latitude:units = "deg" ;
		latitude:missing_value = -1.e+030f ;
	float view_zenith(matchup, nj, ni) ;
		view_zenith:units = "deg" ;
		view_zenith:missing_value = -1.e+030f ;
	float sun_zenith(matchup, nj, ni) ;
		sun_zenith:units = "deg" ;
		sun_zenith:missing_value = -1.e+030f ;
	float delta_azimuth(matchup, nj, ni) ;
		delta_azimuth:units = "deg" ;
		delta_azimuth:missing_value = -1.e+030f ;
	float reflec_1(matchup, nj, ni) ;
		reflec_1:units = "%" ;
		reflec_1:missing_value = -1.e+030f ;
	float reflec_2(matchup, nj, ni) ;
		reflec_2:units = "%" ;
		reflec_2:missing_value = -1.e+030f ;
	float reflec_3a(matchup, nj, ni) ;
		reflec_3a:units = "%" ;
		reflec_3a:missing_value = -1.e+030f ;
	float temp_3b(matchup, nj, ni) ;
		temp_3b:units = "K" ;
		temp_3b:missing_value = -1.e+030f ;
	float temp_4(matchup, nj, ni) ;
		temp_4:units = "K" ;
		temp_4:missing_value = -1.e+030f ;
	float temp_5(matchup, nj, ni) ;
		temp_5:units = "K" ;
		temp_5:missing_value = -1.e+030f ;

// global attributes:
		:title = "AVHRR matchup" ;
		:source = "Version 1.0 of GBCS cloud screening code, IAES, University of Edinburgh, 2011" ;
		:GBCS_rev = "$Rev: 882 $" ;
}
