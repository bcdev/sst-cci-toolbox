netcdf l2p {
dimensions:
    ni = 512 ;
    nj = 40000 ;
    time = 1 ;
variables:
    float lat(nj, ni) ;
        lat:units = "degrees_north" ;
        lat:long_name = "Latitude coordinates" ;
        lat:standard_name = "latitude" ;
        lat:valid_min = -90.0f ;
        lat:valid_max = 90.0f ;
        lat:reference_datum = "geographical coordinates, WGS84 projection" ;
    float lon(nj, ni) ;
        lon:units = "degrees_east" ;
        lon:long_name = "Longitude coordinates" ;
        lon:standard_name = "longitude" ;
        lon:valid_min = -180.0f ;
        lon:valid_max = 180.0f ;
        lon:reference_datum = "geographical coordinates, WGS84 projection" ;
    int time(time) ;
        time:units = "seconds since 1981-01-01 00:00:00" ;
        time:long_name = "reference time of sst file" ;
        time:standard_name = "time" ;
        time:calendar = "gregorian" ;
    short sea_surface_temperature(time, nj, ni) ;
        sea_surface_temperature:_FillValue = -32768s ;
        sea_surface_temperature:units = "kelvin" ;
        sea_surface_temperature:scale_factor = 0.01f ;
        sea_surface_temperature:add_offset = 273.15f ;
        sea_surface_temperature:long_name = "sea surface skin temperature" ;
        sea_surface_temperature:valid_min = -200s;
        sea_surface_temperature:valid_max = 5000s;
        sea_surface_temperature:standard_name = "sea_surface_skin_temperature" ;
        sea_surface_temperature:comment = "Temperature of the skin of the ocean; total uncertainty = sqrt(large_scale_correlated_uncertainty^2 + synoptically_correlated _uncertainty^2 + uncorrelated_uncertainty^2)" ;
        sea_surface_temperature:source = "TBD" ;
        sea_surface_temperature:references = "TBD" ;
        sea_surface_temperature:depth = "10 micrometres" ;
        sea_surface_temperature:coordinates = "lon lat" ;
    short sst_dtime(time, nj, ni) ;
        sst_dtime:_FillValue = -32768s ;
        sst_dtime:units = "seconds" ;
        sst_dtime:long_name = "time difference from reference time" ;
        sst_dtime:valid_min = -32767s ;
        sst_dtime:valid_max = 32767s ;
        sst_dtime:comment = "time plus sst_dtime gives seconds after 1981-01-01 00:00:00" ;
        sst_dtime:coordinates = "lon lat" ;
    byte sses_bias(time, nj, ni) ;
        sses_bias:_FillValue = -128b ;
        sses_bias:units = "kelvin" ;
        sses_bias:scale_factor = 0.01f ;
        sses_bias:add_offset = 0.0f ;
        sses_bias:long_name = "SSES bias factor" ;
        sses_bias:valid_min = -127b ;
        sses_bias:valid_max = 127b ;
        sses_bias:comment = "No SSES biases and standard deviations are available for these data; see large_scale_correlated_uncertainty, synoptically_correlated_uncertainty, uncorrelated_uncertainty adjustment_uncertainty instead" ;
        sses_bias:coordinates = "lon lat" ;
    byte sses_standard_deviation(time, nj, ni) ;
        sses_standard_deviation:_FillValue = -128b ;
        sses_standard_deviation:units = "kelvin" ;
        sses_standard_deviation:scale_factor = 0.01f ;
        sses_standard_deviation:add_offset = 0.0f ;
        sses_standard_deviation:long_name = "SSES standard deviation" ;
        sses_standard_deviation:valid_min = -127b ;
        sses_standard_deviation:valid_max = 127b ;
        sses_standard_deviation:comment = "No SSES biases and standard deviations are available for these data; see large_scale_correlated_uncertainty, synoptically_correlated_uncertainty, uncorrelated_uncertainty adjustment_uncertainty instead" ;
        sses_standard_deviation:coordinates = "lon lat" ;
    short l2p_flags(time, nj, ni) ;
        l2p_flags:long_name = "L2P flags" ;
        l2p_flags:flag_meanings = "microwave land ice lake river spare views channels" ;
        l2p_flags:flag_masks = 1s, 2s, 4s, 8s, 16s, 32s, 64s, 128s ;
        l2p_flags:comment = "These flags are important to use the data" ;
        l2p_flags:coordinates = "lon lat" ;
    byte quality_level(time, nj, ni) ;
        quality_level:long_name = "Quality level of SST pixel" ;
        quality_level:flag_meanings = "no_data bad_data worst_quality low_quality acceptable_quality best_quality" ;
        quality_level:flag_values = 0b, 1b, 2, 3b, 4b, 5b ;
        quality_level:comment = "These are the overall quality indicators and are those used for all GHRSST SSTs" ;
        quality_level:coordinates = "lon lat" ;
    byte wind_speed(time, nj, ni) ;
        wind_speed:_FillValue = -128b ;
        wind_speed:units = "m s-1" ;
        wind_speed:scale_factor = 0.1f ;
        wind_speed:add_offset = 12.7f ;
        wind_speed:long_name = "10m wind speed" ;
        wind_speed:valid_min = -127b ;
        wind_speed:valid_max = 127b ;
        wind_speed:standard_name = "wind_speed" ;
        wind_speed:comment = "Wind speeds sourced from ECMWF ERA Interim reanalysis; wind speeds greater than 25.4 m s-1 are set to 25.4" ;
        wind_speed:coordinates = "lon lat" ;
        wind_speed:height = "10 m" ;
        wind_speed:source = "TBD" ;
        wind_speed:references = "TBD" ;
        wind_speed:time_offset = 0b ;
    short tos(time, nj, ni) ;
        tos:_FillValue = -32768s ;
        tos:units = "kelvin" ;
        tos:scale_factor = 0.01f ;
        tos:add_offset = 273.15f ;
        tos:long_name = "sea surface temperature at 0.2 m" ;
        tos:valid_min = -200s ;
        tos:valid_max = 5000s ;
        tos:standard_name = "sea_water_temperature" ;
        tos:comment = "Temperature of the ocean at 20 cm depth; total uncertainty = sqrt(large_scale_correlated_uncertainty^2 + synoptically_correlated_uncertainty^2 + uncorrelated_uncertainty^2 + adjustment_uncertainty^2)" ;
        tos:coordinates = "lon lat" ;
        tos:depth = "0.2 m" ;
        tos:source = "TBD" ;
        tos:references = "TBD" ;
    short large_scale_correlated_uncertainty(time, nj, ni) ;
        large_scale_correlated_uncertainty:_FillValue = -32768s ;
        large_scale_correlated_uncertainty:units = "kelvin" ;
        large_scale_correlated_uncertainty:scale_factor = 0.01f ;
        large_scale_correlated_uncertainty:add_offset = 0.0f ;
        large_scale_correlated_uncertainty:long_name = "Uncertainty from errors likely to be correlated over large scales" ;
        large_scale_correlated_uncertainty:valid_min = 0s ;
        large_scale_correlated_uncertainty:valid_max = 5000s ;
        large_scale_correlated_uncertainty:comment = "Component of uncertainty that is correlated over large scales; can be combined with other uncertainty estimates to form a total uncertainty" ;
        large_scale_correlated_uncertainty:coordinates = "lon lat" ;
        large_scale_correlated_uncertainty:references = "TBD" ;
    short synoptically_correlated_uncertainty(time, nj, ni) ;
        synoptically_correlated_uncertainty:_FillValue = -32768s ;
        synoptically_correlated_uncertainty:units = "kelvin" ;
        synoptically_correlated_uncertainty:scale_factor = 0.01f ;
        synoptically_correlated_uncertainty:add_offset = 0.0f ;
        synoptically_correlated_uncertainty:long_name = "Uncertainty from errors likely to be correlated over synoptic scales" ;
        synoptically_correlated_uncertainty:valid_min = 0s ;
        synoptically_correlated_uncertainty:valid_max = 5000s ;
        synoptically_correlated_uncertainty:comment = "Component of uncertainty that is correlated over synoptic scales; can be combined with other uncertainty estimates to form a total uncertainty" ;
        synoptically_correlated_uncertainty:coordinates = "lon lat" ;
        synoptically_correlated_uncertainty:references = "TBD" ;
        synoptically_correlated_uncertainty:correlation_length_scale = "100 km" ;
        synoptically_correlated_uncertainty:correlation_time_scale = "1 day" ;
    short uncorrelated_uncertainty(time, nj, ni) ;
        uncorrelated_uncertainty:_FillValue = -32768s ;
        uncorrelated_uncertainty:units = "kelvin" ;
        uncorrelated_uncertainty:scale_factor = 0.01f ;
        uncorrelated_uncertainty:add_offset = 0.0f ;
        uncorrelated_uncertainty:long_name = "Uncertainty from errors likely to be uncorrelated between SSTs" ;
        uncorrelated_uncertainty:valid_min = 0s ;
        uncorrelated_uncertainty:valid_max = 5000s ;
        uncorrelated_uncertainty:comment = "Component of uncertainty that is uncorrelated between SSTs; can be combined with other uncertainty estimates to form a total uncertainty" ;
        uncorrelated_uncertainty:coordinates = "lon lat" ;
        uncorrelated_uncertainty:references = "TBD" ;
    short adjustment_uncertainty(time, nj, ni) ;
        adjustment_uncertainty:_FillValue = -32768s ;
        adjustment_uncertainty:units = "kelvin" ;
        adjustment_uncertainty:scale_factor = 0.01f ;
        adjustment_uncertainty:add_offset = 0.0f ;
        adjustment_uncertainty:long_name = "Time and depth adjustment uncertainty" ;
        adjustment_uncertainty:valid_min = 0s ;
        adjustment_uncertainty:valid_max = 5000s ;
        adjustment_uncertainty:comment = "Adjustment uncertainty; can be combined with other uncertainty estimates to form a total uncertainty" ;
        adjustment_uncertainty:coordinates = "lon lat" ;
        adjustment_uncertainty:references = "TBD" ;

// global attributes:
        :Conventions = "CF-1.4" ;
        :title = "ESA SST CCI AATSR L2P product" ;
        :summary = "AATSR L2P product from the ESA SST CCI project, produced using <algorithm name>" ;
        :references = "TBD" ;
        :institution = "ESACCI" ;
        :history = "" ;
        :license = "GHRSST protocol describes data use as free and open" ;
        :id = "TBD" ;
        :naming_authority = "org.ghrsst" ;
        :product_version = "TBD" ;
        :uuid = "TBD" ;
        :gds_version_id = "2.0" ;
        :netcdf_version_id = "4.1.3" ;
        :date_created = "20120131T120000Z" ;
        :file_quality_level = 0 ;
        :spatial_resolution = "1 km" ;
        :start_time = "20120131070000Z" ;
        :time_coverage_start = "20120131070000Z" ;
        :stop_time = "20120131083000Z" ;
        :source = "AATSR-ESA-L1-v2.0" ;
        :platform = "Envisat" ;
        :sensor = "AATSR" ;
        :metadata_conventions = "Unidata Dataset Discovery v1.0" ;
        :metadata_link = "TBD" ;
        :keywords = "Oceans > Ocean > Temperature > Sea Surface Temperature" ;
        :keywords_vocabulary = "NASA Global Change Master Directory (GCMD) Science Keywords" ;
        :standard_name_vocabulary = "NetCDF Climate and Forecast (CF) Metadata Convention" ;
        :geospatial_lat_units = "degrees_north" ;
        :geospatial_lon_units = "degrees_east" ;
        :acknowledgment = "Funded by ESA" ;
        :creator_name = "ESA SST CCI" ;
        :creator_email = "science.lead er@esa-sst- cci.org" ;
        :creator_url = "http://www.es a-sst-cci.org/" ;
        :project = "European Space Agency Sea Surface Temperature Climate Change Initiative" ;
        :publisher_name = "The GHRSST Project Office" ;
        :publisher_email = "ghrsst- po@nceo.ac.uk" ;
        :publisher_url = "http://www.g hrsst.org" ;
        :comment = "These data were produced at ESACCI as part of the ESA SST CCI project. This file does not include single sensor error statistics. Alternative uncertainty statistics are provided instead. See the comment attributes to the sea_surface temperature and tos variables for information about uncertainty estimates" ;
        :northernmost_latitude = 90.0f ;
        :southernmost_latitude = -90.0f ;
        :easternmost_longitude = 180.0f ;
        :westernmost_longitude = -180.0f ;
        :processing_level = "L2P" ;
        :cdm_data_type = "swath" ;
}