netcdf arc3_output_mmd {
dimensions:
	ni = 101 ;
	nj = 101 ;
	record = UNLIMITED ; // (169 currently)
	depth = 3 ;
variables:
	int matchup_id(record) ;
	float lon(record, nj, ni) ;
		lon:long_name = "Longitude coordinates" ;
		lon:standard_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:valid_min = -180.f ;
		lon:valid_max = 180.f ;
	float lat(record, nj, ni) ;
		lat:long_name = "Latitude coordinates" ;
		lat:standard_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:valid_min = -90.f ;
		lat:valid_max = 90.f ;
	float atsr.3.cloud_mask.bayes_nadir_min(record, nj, ni) ;
		atsr.3.cloud_mask.bayes_nadir_min:long_name = "Probability of clear-sky" ;
		atsr.3.cloud_mask.bayes_nadir_min:_FillValue = -999.f ;
		atsr.3.cloud_mask.bayes_nadir_min:valid_min = 0.f ;
		atsr.3.cloud_mask.bayes_nadir_min:valid_max = 1.f ;
	float atsr.3.cloud_mask.bayes_dual_max(record, nj, ni) ;
		atsr.3.cloud_mask.bayes_dual_max:long_name = "Probability of clear-sky" ;
		atsr.3.cloud_mask.bayes_dual_max:_FillValue = -999.f ;
		atsr.3.cloud_mask.bayes_dual_max:valid_min = 0.f ;
		atsr.3.cloud_mask.bayes_dual_max:valid_max = 1.f ;
	short atsr.3.sea_surface_temperature.ARC.N2(record, nj, ni) ;
		atsr.3.sea_surface_temperature.ARC.N2:standard_name = "sea_surface_skin_temperature" ;
		atsr.3.sea_surface_temperature.ARC.N2:long_name = "sea surface skin temperature" ;
		atsr.3.sea_surface_temperature.ARC.N2:units = "kelvin" ;
		atsr.3.sea_surface_temperature.ARC.N2:_FillValue = -32768s ;
		atsr.3.sea_surface_temperature.ARC.N2:scale_factor = 0.01f ;
		atsr.3.sea_surface_temperature.ARC.N2:add_offset = 273.15f ;
		atsr.3.sea_surface_temperature.ARC.N2:valid_min = -200s ;
		atsr.3.sea_surface_temperature.ARC.N2:valid_max = 5000s ;
	short atsr.3.sea_surface_temperature.op.N2(record, nj, ni) ;
		atsr.3.sea_surface_temperature.op.N2:standard_name = "sea_surface_skin_temperature" ;
		atsr.3.sea_surface_temperature.op.N2:long_name = "sea surface skin temperature" ;
		atsr.3.sea_surface_temperature.op.N2:units = "kelvin" ;
		atsr.3.sea_surface_temperature.op.N2:_FillValue = -32768s ;
		atsr.3.sea_surface_temperature.op.N2:scale_factor = 0.01f ;
		atsr.3.sea_surface_temperature.op.N2:add_offset = 273.15f ;
		atsr.3.sea_surface_temperature.op.N2:valid_min = -200s ;
		atsr.3.sea_surface_temperature.op.N2:valid_max = 5000s ;
	float atsr.3.saharan_dust_index.2(record, nj, ni) ;
		atsr.3.saharan_dust_index.2:standard_name = "ASDI2" ;
		atsr.3.saharan_dust_index.2:long_name = "ATSR Saharan Dust Index from 2 channel algorithm" ;
		atsr.3.saharan_dust_index.2:units = "kelvin" ;

// global attributes:
		:netcdf_version_id = "\"3.6.3\" of Jul 30 2008 18:07:43 $" ;
		:date_created = "20110411T161448Z" ;
		:history = "Created using GBCS library $Rev: 1215 $" ;
		:Conventions = "CF-1.4, Unidata Observation Dataset v1.0" ;
		:institution = "ESACCI" ;
		:comment = "These data were produced at University of Edinburgh as part of the ESA SST CCI project." ;
		:licence = "GHRSST protocol describes data use as free and open." ;
		:product_version = "0.1" ;
		:gds_version_id = "2.0" ;
		:metadata_conventions = "Unidata Dataset Discovery v1.0" ;
		:keywords = "Oceans > Ocean Temperature > Sea Surface Temperature" ;
		:keywords_vocabulary = "NASA Global change Master Directory (GCMD) Science Keywords" ;
		:standard_name_vocabulary = "NetCDF Climate and Forecast (CF) Metadata Convention" ;
		:acknowledgment = "Funded by ESA" ;
		:creator_name = "ESA SST CCI" ;
		:creator_email = "science.leader@esa-sst-cci.org" ;
		:creator_url = "http://www.esa-sst-cci.org/" ;
		:project = "European Space Agency Sea Surface Temperature Climate Change Initiative" ;
		:publisher_name = "The GHRSST Project Office" ;
		:publisher_url = "http://www.ghrsst.org" ;
		:publisher_email = "ghrsst-po@nceo.ac.uk" ;
}
